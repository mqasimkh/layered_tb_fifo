class env;
endclass: env